module tokenizer

// token:=['\n', 'for', ' ', 'i', ',', 'char', ' ', 'in', ' ', 'enumerate', '(', 'str', 'in', 'g', ')', ':', '\n', ' ', ' ', ' ', ' ', 'if', ' ', 'char', ' ', '!', '=', ' ', 'white_space', ':', '\n', '         ', '#', ' ', 'adding', ' ', 'a', ' ', 'char', ' ', 'each', ' ', 'time', '\n', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', 'lexeme', ' ', '+', '=', ' ', 'char', ' ', '\n', ' ', ' ', ' ', ' ', '#', 'print', '(', 'lexeme', ')', '\n', '    ', '#', ' ', 'prevents', ' ', 'error', '\n', ' ', ' ', ' ', ' ', 'if', ' ', 'i', '+', '1', ' ', '<', ' ', 'len', '(', 'str', 'in', 'g', ')', ':', '\n', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', 'if', ' ', 'str', 'in', 'g', '[', 'i', '+', '1', ']', ' ', '=', '=', ' ', 'white_space', ' ', 'or', ' ', 'str', 'in', 'g', '[', 'i', '+', '1', ']', ' ', 'in', ' ', 'KEYWORDS', ' ', 'or', ' ', 'lexeme', ' ', 'in', ' ', 'KEYWORDS', ':', ' ', '#', ' ', 'if', ' ', 'next', ' ', 'char', ' ', '=', '=', ' ', ''', ' ', ''', '\n', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', 'if', ' ', 'lexeme', ' ', '!', '=', ' ', ''', ''', ':', '\n', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', 'a', '.', 'append', '(', 'lexeme', '.', 'replace', '(', ''', '\n', ''', ',', ' ', ''', '<', 'newline', '>', ''', ')', ')', '\n', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', 'print', '(', 'lexeme', '.', 'replace', '(', ''', '\n', ''', ',', ' ', ''', '<', 'newline', '>', ''', ')', ')', '\n', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', ' ', 'lexeme', ' ', '=', ' ', ''', ''', '\n', 'print', '(', 'a', ')', '\n']