module parser

// Original author : Saptak Bhoumik
fn factor() {
}

fn term() {
}

fn expression() {
}
