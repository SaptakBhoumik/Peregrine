module parser
// Original author : Saptak Bhoumik
// enum Num{}
fn factor(){
	// mut value := 0
    // if (token == '(') {
    //     match('(')
    //     	value = expr()
    //     match(')')
    // } else {
    //     value = token_val
    //     match(Num)
    // }
    // return value
}
fn term(){

}
fn expression(){

}