module tokenizer

// lis = [" ","1","f","2"," " ,"3", "world", "hello", "hel", "ho", "hlo"]

// count = 0

// for i in lis:
//     count += 1
//     if i == " ":
//         break

// lis[count] = lis[count] + "".join([str(x) for x in lis[count + 1 : len(lis)]]) 

// lis = "".join(str(lis[0:count + 1])).replace("'", "").replace(",", " ").replace("[", "").replace("]", "")

// print(lis.split())